`define SOC_SPI1_BASE_ADDRESS 32'h20000200
`define SOC_SPI1_END_ADDRESS 32'h2000027F

`define SOC_SPI2_BASE_ADDRESS 32'h20000280
`define SOC_SPI2_END_ADDRESS 32'h200002FF
`define OFFSET 4
