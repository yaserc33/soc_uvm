package common_pkg;

typedef enum logic[0:0] {
	FALSE,
	TRUE
} onebit_sig_e;

endpackage