package soc_pkg ; 
 `include "uvm_macros.svh"
 import uvm_pkg::*;
 import spi_pkg::*;
 import wb_pkg::*;
import clock_and_reset_pkg::*;
import spi_module_pkg::*;


// import uart_pkg::*;
// import wb_pkg::*;

`include "wb_ref_model.sv"
`include "soc_scb.sv"
`include "soc_ref_env.sv"



endpackage